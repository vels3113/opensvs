* y.spice
M1 Vout Vin VDD VDD PMOS w=800n l=400n
M2 Vout Vin VDD VDD PMOS w=800n l=400n
M3 Vout Vin 0 0 NMOS w=800n l=400n