* SPICE3 file created from map9v3.ext - technology: scmos

.subckt BUFX2 Y gnd A vdd
M1000 vdd A a_10_30# vdd pfet w=4u l=0.4u
+ ad=8.8p pd=18.4u as=4p ps=10u 
M1001 Y a_10_30# vdd vdd pfet w=8u l=0.4u
+ ad=8p pd=18u as=0p ps=0u 
M1002 gnd A a_10_30# Gnd nfet w=2u l=0.4u
+ ad=4.4p pd=10.4u as=2p ps=6u 
M1003 Y a_10_30# gnd Gnd nfet w=4u l=0.4u
+ ad=4p pd=10u as=0p ps=0u 
.ends

.subckt DFFPOSX1 gnd CLK D Q vdd
M1000 vdd CLK a_10_30# vdd pfet w=8u l=0.4u
+ ad=26p pd=57.2u as=8p ps=18u 
M1001 a_85_370# D vdd vdd pfet w=4u l=0.4u
+ ad=3.2p pd=9.6u as=0p ps=0u 
M1002 a_110_30# CLK a_85_370# vdd pfet w=4u l=0.4u
+ ad=4.8p pd=10.4u as=0p ps=0u 
M1003 a_155_370# a_10_30# a_110_30# vdd pfet w=4u l=0.4u
+ ad=3.2p pd=9.6u as=0p ps=0u 
M1004 vdd a_170_20# a_155_370# vdd pfet w=4u l=0.4u
+ ad=0p pd=0u as=0p ps=0u 
M1005 a_170_20# a_110_30# vdd vdd pfet w=4u l=0.4u
+ ad=4p pd=10u as=0p ps=0u 
M1006 a_305_370# a_170_20# vdd vdd pfet w=4u l=0.4u
+ ad=2.4p pd=9.2u as=0p ps=0u 
M1007 a_330_30# a_10_30# a_305_370# vdd pfet w=4u l=0.4u
+ ad=6p pd=11.2u as=0p ps=0u 
M1008 a_380_420# CLK a_330_30# vdd pfet w=2u l=0.4u
+ ad=1.2p pd=5.2u as=0p ps=0u 
M1009 vdd Q a_380_420# vdd pfet w=2u l=0.4u
+ ad=0p pd=0u as=0p ps=0u 
M1010 gnd CLK a_10_30# Gnd nfet w=4u l=0.4u
+ ad=13.6p pd=33.6u as=4p ps=10u 
M1011 Q a_330_30# vdd vdd pfet w=8u l=0.4u
+ ad=8p pd=18u as=0p ps=0u 
M1012 a_85_30# D gnd Gnd nfet w=2u l=0.4u
+ ad=1.2p pd=5.2u as=0p ps=0u 
M1013 a_110_30# a_10_30# a_85_30# Gnd nfet w=2u l=0.4u
+ ad=2.8p pd=6.8u as=0p ps=0u 
M1014 a_155_30# CLK a_110_30# Gnd nfet w=2u l=0.4u
+ ad=1.2p pd=5.2u as=0p ps=0u 
M1015 gnd a_170_20# a_155_30# Gnd nfet w=2u l=0.4u
+ ad=0p pd=0u as=0p ps=0u 
M1016 a_170_20# a_110_30# gnd Gnd nfet w=2u l=0.4u
+ ad=2p pd=6u as=0p ps=0u 
M1017 a_305_30# a_170_20# gnd Gnd nfet w=2u l=0.4u
+ ad=1.2p pd=5.2u as=0p ps=0u 
M1018 a_330_30# CLK a_305_30# Gnd nfet w=2u l=0.4u
+ ad=3.2p pd=7.2u as=0p ps=0u 
M1019 a_380_30# a_10_30# a_330_30# Gnd nfet w=2u l=0.4u
+ ad=1.2p pd=5.2u as=0p ps=0u 
M1020 gnd Q a_380_30# Gnd nfet w=2u l=0.4u
+ ad=0p pd=0u as=0p ps=0u 
M1021 Q a_330_30# gnd Gnd nfet w=4u l=0.4u
+ ad=4p pd=10u as=0p ps=0u 
.ends

.subckt INVX1 Y gnd A vdd
M1000 Y A vdd vdd pfet w=4u l=0.4u
+ ad=4p pd=10u as=4p ps=10u 
M1001 Y A gnd Gnd nfet w=2u l=0.4u
+ ad=2p pd=6u as=2p ps=6u 
.ends

.subckt NAND2X1 Y gnd A B vdd
M1000 Y A vdd vdd pfet w=4u l=0.4u
+ ad=4.8p pd=10.4u as=8p ps=20u 
M1001 vdd B Y vdd pfet w=4u l=0.4u
+ ad=0p pd=0u as=0p ps=0u 
M1002 a_45_30# A gnd Gnd nfet w=4u l=0.4u
+ ad=2.4p pd=9.2u as=4p ps=10u 
M1003 Y B a_45_30# Gnd nfet w=4u l=0.4u
+ ad=4p pd=10u as=0p ps=0u 
.ends

.subckt OAI21X1 Y gnd A B C vdd
M1000 a_45_270# A vdd vdd pfet w=8u l=0.4u
+ ad=4.8p pd=17.2u as=12p ps=28u 
M1001 Y B a_45_270# vdd pfet w=8u l=0.4u
+ ad=8.8p pd=18.4u as=0p ps=0u 
M1002 vdd C Y vdd pfet w=4u l=0.4u
+ ad=0p pd=0u as=0p ps=0u 
M1003 gnd A a_10_30# Gnd nfet w=4u l=0.4u
+ ad=4.8p pd=10.4u as=8.8p ps=20.4u 
M1004 a_10_30# B gnd Gnd nfet w=4u l=0.4u
+ ad=0p pd=0u as=0p ps=0u 
M1005 Y C a_10_30# Gnd nfet w=4u l=0.4u
+ ad=4p pd=10u as=0p ps=0u 
.ends

.subckt AOI21X1 Y gnd A B C vdd
M1000 vdd A a_10_270# vdd pfet w=8u l=0.4u
+ ad=9.6p pd=18.4u as=17.6p ps=36.4u 
M1001 a_10_270# B vdd vdd pfet w=8u l=0.4u
+ ad=0p pd=0u as=0p ps=0u 
M1002 Y C a_10_270# vdd pfet w=8u l=0.4u
+ ad=8p pd=18u as=0p ps=0u 
M1003 a_60_30# A gnd Gnd nfet w=4u l=0.4u
+ ad=2.4p pd=9.2u as=6p ps=16u 
M1004 Y B a_60_30# Gnd nfet w=4u l=0.4u
+ ad=4.4p pd=10.4u as=0p ps=0u 
M1005 gnd C Y Gnd nfet w=2u l=0.4u
+ ad=0p pd=0u as=0p ps=0u 
.ends

.subckt OAI22X1 Y gnd A B C D vdd
M1000 a_45_270# A vdd vdd pfet w=8u l=0.4u
+ ad=4.8p pd=17.2u as=16p ps=36u 
M1001 Y B a_45_270# vdd pfet w=8u l=0.4u
+ ad=19.2p pd=20.8u as=0p ps=0u 
M1002 a_140_270# D Y vdd pfet w=8u l=0.4u
+ ad=4.8p pd=17.2u as=0p ps=0u 
M1003 vdd C a_140_270# vdd pfet w=8u l=0.4u
+ ad=0p pd=0u as=0p ps=0u 
M1004 gnd A a_10_30# Gnd nfet w=4u l=0.4u
+ ad=4.8p pd=10.4u as=12.8p ps=30.4u 
M1005 a_10_30# B gnd Gnd nfet w=4u l=0.4u
+ ad=0p pd=0u as=0p ps=0u 
M1006 Y D a_10_30# Gnd nfet w=4u l=0.4u
+ ad=4.8p pd=10.4u as=0p ps=0u 
M1007 a_10_30# C Y Gnd nfet w=4u l=0.4u
+ ad=0p pd=0u as=0p ps=0u 
.ends

.subckt MUX2X1 Y gnd B A vdd S
M1000 vdd S a_10_50# vdd pfet w=4u l=0.4u
+ ad=16.32p pd=36.4u as=4p ps=10u 
M1001 a_85_250# B vdd vdd pfet w=8u l=0.4u
+ ad=4.8p pd=17.2u as=0p ps=0u 
M1002 Y S a_85_250# vdd pfet w=8u l=0.4u
+ ad=9.92p pd=20u as=0p ps=0u 
M1003 a_150_270# a_10_50# Y vdd pfet w=8u l=0.4u
+ ad=4.8p pd=17.2u as=0p ps=0u 
M1004 vdd A a_150_270# vdd pfet w=8u l=0.4u
+ ad=0p pd=0u as=0p ps=0u 
M1005 gnd S a_10_50# Gnd nfet w=2u l=0.4u
+ ad=8.24p pd=20.4u as=2p ps=6u 
M1006 a_85_50# B gnd Gnd nfet w=4u l=0.4u
+ ad=2.4p pd=9.2u as=0p ps=0u 
M1007 Y a_10_50# a_85_50# Gnd nfet w=4u l=0.4u
+ ad=4.8p pd=10.4u as=0p ps=0u 
M1008 a_150_50# S Y Gnd nfet w=4u l=0.4u
+ ad=2.4p pd=9.2u as=0p ps=0u 
M1009 gnd A a_150_50# Gnd nfet w=4u l=0.4u
+ ad=0p pd=0u as=0p ps=0u 
.ends

.subckt AOI22X1 Y gnd A B C D vdd
M1000 vdd A a_10_270# vdd pfet w=8u l=0.4u
+ ad=9.6p pd=18.4u as=25.6p ps=54.4u 
M1001 a_10_270# B vdd vdd pfet w=8u l=0.4u
+ ad=0p pd=0u as=0p ps=0u 
M1002 Y D a_10_270# vdd pfet w=8u l=0.4u
+ ad=9.6p pd=18.4u as=0p ps=0u 
M1003 a_10_270# C Y vdd pfet w=8u l=0.4u
+ ad=0p pd=0u as=0p ps=0u 
M1004 a_55_30# A gnd Gnd nfet w=4u l=0.4u
+ ad=2.4p pd=9.2u as=8p ps=20u 
M1005 Y B a_55_30# Gnd nfet w=4u l=0.4u
+ ad=8p pd=12u as=0p ps=0u 
M1006 a_140_30# D Y Gnd nfet w=4u l=0.4u
+ ad=2.4p pd=9.2u as=0p ps=0u 
M1007 gnd C a_140_30# Gnd nfet w=4u l=0.4u
+ ad=0p pd=0u as=0p ps=0u 
.ends

.subckt OR2X1 Y gnd A B vdd
M1000 a_45_270# A a_10_270# vdd pfet w=8u l=0.4u
+ ad=4.8p pd=17.2u as=8p ps=18u 
M1001 vdd B a_45_270# vdd pfet w=8u l=0.4u
+ ad=8.8p pd=18.4u as=0p ps=0u 
M1002 Y a_10_270# vdd vdd pfet w=4u l=0.4u
+ ad=4p pd=10u as=0p ps=0u 
M1003 a_10_270# A gnd Gnd nfet w=2u l=0.4u
+ ad=2.4p pd=6.4u as=4.4p ps=12.4u 
M1004 gnd B a_10_270# Gnd nfet w=2u l=0.4u
+ ad=0p pd=0u as=0p ps=0u 
M1005 Y a_10_270# gnd Gnd nfet w=2u l=0.4u
+ ad=2p pd=6u as=0p ps=0u 
.ends

.subckt NAND3X1 Y gnd A B C vdd
M1000 Y A vdd vdd pfet w=4u l=0.4u
+ ad=8.8p pd=20.4u as=8.8p ps=20.4u 
M1001 vdd B Y vdd pfet w=4u l=0.4u
+ ad=0p pd=0u as=0p ps=0u 
M1002 Y C vdd vdd pfet w=4u l=0.4u
+ ad=0p pd=0u as=0p ps=0u 
M1003 a_45_30# A gnd Gnd nfet w=6u l=0.4u
+ ad=3.6p pd=13.2u as=6p ps=14u 
M1004 a_70_30# B a_45_30# Gnd nfet w=6u l=0.4u
+ ad=3.6p pd=13.2u as=0p ps=0u 
M1005 Y C a_70_30# Gnd nfet w=6u l=0.4u
+ ad=6p pd=14u as=0p ps=0u 
.ends

.subckt NOR2X1 Y gnd A B vdd
M1000 a_45_270# A vdd vdd pfet w=8u l=0.4u
+ ad=4.8p pd=17.2u as=8p ps=18u 
M1001 Y B a_45_270# vdd pfet w=8u l=0.4u
+ ad=8p pd=18u as=0p ps=0u 
M1002 Y A gnd Gnd nfet w=2u l=0.4u
+ ad=2.4p pd=6.4u as=4p ps=12u 
M1003 gnd B Y Gnd nfet w=2u l=0.4u
+ ad=0p pd=0u as=0p ps=0u 
.ends


* Top level circuit map9v3

X0 dp<8> INVX1_3/gnd BUFX2_10/A INVX1_3/vdd BUFX2
X1 INVX1_3/gnd clock OAI21X1_19/Y BUFX2_10/A INVX1_3/vdd DFFPOSX1
X2 INVX1_6/Y INVX1_3/gnd INVX1_6/A INVX1_3/vdd INVX1
X3 OAI21X1_19/C INVX1_3/gnd OR2X1_2/Y BUFX2_10/A INVX1_3/vdd NAND2X1
X4 OAI21X1_19/Y INVX1_3/gnd OR2X1_3/Y MUX2X1_1/A OAI21X1_19/C INVX1_3/vdd OAI21X1
X5 NAND2X1_20/Y INVX1_3/gnd OR2X1_2/Y BUFX2_4/A INVX1_3/vdd NAND2X1
X6 INVX1_3/gnd clock OAI21X1_3/Y BUFX2_9/A INVX1_3/vdd DFFPOSX1
X7 OAI21X1_3/Y INVX1_3/gnd INVX1_9/Y OR2X1_3/Y NAND2X1_3/Y INVX1_3/vdd OAI21X1
X8 NAND2X1_3/Y INVX1_3/gnd OR2X1_2/Y BUFX2_9/A INVX1_3/vdd NAND2X1
X9 dp<6> INVX1_3/gnd BUFX2_9/A INVX1_3/vdd BUFX2
X10 INVX1_3/gnd clock OAI21X1_18/Y BUFX2_3/A INVX1_3/vdd DFFPOSX1
X11 dp<5> INVX1_3/gnd BUFX2_3/A INVX1_3/vdd BUFX2
X12 OAI21X1_18/Y INVX1_3/gnd OR2X1_3/Y INVX1_10/Y NAND2X1_22/Y INVX1_3/vdd OAI21X1
X13 NAND2X1_22/Y INVX1_3/gnd OR2X1_2/Y BUFX2_3/A INVX1_3/vdd NAND2X1
X14 INVX1_3/gnd clock OAI22X1_3/Y INVX1_9/A INVX1_3/vdd DFFPOSX1
X15 INVX1_3/gnd clock OR2X1_2/B BUFX2_5/A INVX1_3/vdd DFFPOSX1
X16 done INVX1_3/gnd BUFX2_5/A INVX1_3/vdd BUFX2
X17 INVX1_3/gnd clock INVX1_1/Y OR2X1_2/B INVX1_3/vdd DFFPOSX1
X18 INVX1_3/gnd clock reset AOI21X1_1/C INVX1_3/vdd DFFPOSX1
X19 AOI21X1_1/Y INVX1_3/gnd INVX1_3/Y start AOI21X1_1/C INVX1_3/vdd AOI21X1
X20 INVX1_3/gnd clock start INVX1_3/A INVX1_3/vdd DFFPOSX1
X21 INVX1_3/Y INVX1_3/gnd INVX1_3/A INVX1_3/vdd INVX1
X22 dp<7> INVX1_3/gnd BUFX2_4/A INVX1_4/vdd BUFX2
X23 INVX1_3/gnd clock OAI21X1_11/Y BUFX2_4/A INVX1_4/vdd DFFPOSX1
X24 INVX1_29/Y INVX1_3/gnd INVX1_29/A INVX1_4/vdd INVX1
X25 INVX1_3/gnd clock OAI22X1_9/Y INVX1_29/A INVX1_4/vdd DFFPOSX1
X26 OAI21X1_11/Y INVX1_3/gnd OR2X1_3/Y INVX1_29/Y NAND2X1_20/Y INVX1_4/vdd OAI21X1
X27 OAI22X1_9/Y INVX1_3/gnd OAI22X1_3/A INVX1_9/Y OR2X1_1/Y INVX1_29/Y INVX1_4/vdd OAI22X1
X28 OAI22X1_13/Y INVX1_3/gnd OAI22X1_3/A INVX1_29/Y OR2X1_1/Y MUX2X1_1/A INVX1_4/vdd OAI22X1
X29 OAI22X1_3/Y INVX1_3/gnd OAI22X1_3/A INVX1_10/Y OR2X1_1/Y INVX1_9/Y INVX1_4/vdd OAI22X1
X30 INVX1_3/gnd clock OAI22X1_13/Y MUX2X1_1/B INVX1_4/vdd DFFPOSX1
X31 MUX2X1_1/A INVX1_3/gnd MUX2X1_1/B INVX1_4/vdd INVX1
X32 MUX2X1_1/Y INVX1_3/gnd MUX2X1_1/B MUX2X1_1/A INVX1_4/vdd MUX2X1_1/S MUX2X1
X33 MUX2X1_1/S INVX1_3/gnd INVX1_9/Y INVX1_10/Y INVX1_9/A INVX1_10/A INVX1_4/vdd AOI22X1
X34 INVX1_9/Y INVX1_3/gnd INVX1_9/A INVX1_4/vdd INVX1
X35 OR2X1_2/Y INVX1_3/gnd INVX1_1/A OR2X1_2/B INVX1_4/vdd OR2X1
X36 OR2X1_1/Y INVX1_3/gnd reset OR2X1_1/B INVX1_4/vdd OR2X1
X37 INVX1_7/Y INVX1_3/gnd reset INVX1_4/vdd INVX1
X38 OAI21X1_9/C INVX1_3/gnd OAI21X1_9/B INVX1_7/Y INVX1_1/Y INVX1_4/vdd NAND3X1
X39 OAI21X1_9/Y INVX1_3/gnd INVX1_1/Y OAI21X1_9/B OAI21X1_9/C INVX1_4/vdd OAI21X1
X40 INVX1_3/gnd clock OAI21X1_9/Y INVX1_1/A INVX1_4/vdd DFFPOSX1
X41 INVX1_1/Y INVX1_3/gnd INVX1_1/A INVX1_4/vdd INVX1
X42 OR2X1_1/B INVX1_3/gnd reset AOI21X1_1/Y INVX1_1/Y INVX1_4/vdd OAI21X1
X43 INVX1_39/Y INVX1_3/gnd INVX1_39/A INVX1_4/vdd INVX1
X44 INVX1_3/gnd clock INVX1_39/Y OR2X1_6/A INVX1_4/vdd DFFPOSX1
X45 OAI21X1_2/Y INVX1_3/gnd INVX1_4/A INVX1_1/Y INVX1_5/Y INVX1_4/vdd OAI21X1
X46 INVX1_3/gnd clock OAI21X1_2/Y INVX1_4/A INVX1_4/vdd DFFPOSX1
X47 dp<2> INVX1_4/gnd BUFX2_7/A INVX1_4/vdd BUFX2
X48 INVX1_4/gnd clock OAI21X1_14/Y BUFX2_7/A INVX1_4/vdd DFFPOSX1
X49 OAI21X1_14/C INVX1_4/gnd OR2X1_2/Y BUFX2_7/A INVX1_4/vdd NAND2X1
X50 OAI21X1_14/Y INVX1_4/gnd INVX1_6/Y OR2X1_3/Y OAI21X1_14/C INVX1_4/vdd OAI21X1
X51 INVX1_4/gnd clock OAI22X1_6/Y INVX1_21/A INVX1_4/vdd DFFPOSX1
X52 INVX1_4/gnd clock OAI22X1_7/Y INVX1_27/A INVX1_4/vdd DFFPOSX1
X53 INVX1_27/Y INVX1_4/gnd INVX1_27/A INVX1_4/vdd INVX1
X54 OAI22X1_11/Y INVX1_4/gnd OAI22X1_3/A INVX1_27/Y OR2X1_1/Y INVX1_10/Y INVX1_4/vdd OAI22X1
X55 INVX1_10/Y INVX1_4/gnd INVX1_10/A INVX1_4/vdd INVX1
X56 INVX1_4/gnd clock INVX1_32/Y INVX1_31/A INVX1_4/vdd DFFPOSX1
X57 INVX1_32/Y INVX1_4/gnd INVX1_32/A INVX1_4/vdd INVX1
X58 INVX1_4/gnd clock INVX1_33/Y INVX1_20/A INVX1_4/vdd DFFPOSX1
X59 OAI22X1_3/A INVX1_4/gnd INVX1_7/Y INVX1_1/A INVX1_4/vdd NAND2X1
X60 INVX1_33/Y INVX1_4/gnd INVX1_33/A INVX1_4/vdd INVX1
X61 INVX1_24/Y INVX1_4/gnd INVX1_24/A INVX1_4/vdd INVX1
X62 OAI21X1_9/B INVX1_4/gnd INVX1_7/Y INVX1_18/A NAND3X1_4/Y INVX1_4/vdd NAND3X1
X63 NAND3X1_4/Y INVX1_4/gnd INVX1_24/Y NOR2X1_3/Y NOR2X1_4/Y INVX1_4/vdd NAND3X1
X64 NOR2X1_4/Y INVX1_4/gnd NOR2X1_4/A NOR2X1_4/B INVX1_4/vdd NOR2X1
X65 INVX1_39/A INVX1_4/gnd INVX1_1/A NOR2X1_4/A AOI21X1_7/C INVX1_4/vdd AOI21X1
X66 NAND2X1_17/Y INVX1_4/gnd OR2X1_6/Y INVX1_20/A INVX1_4/vdd NAND2X1
X67 NOR2X1_4/A INVX1_4/gnd OR2X1_6/Y NAND2X1_15/Y INVX1_4/vdd NAND2X1
X68 NAND2X1_15/Y INVX1_4/gnd OR2X1_6/B OR2X1_6/A INVX1_4/vdd NAND2X1
X69 OR2X1_6/Y INVX1_4/gnd OR2X1_6/A OR2X1_6/B INVX1_4/vdd OR2X1
X70 INVX1_5/A INVX1_4/gnd INVX1_2/Y INVX1_18/A INVX1_4/Y OR2X1_1/B INVX1_4/vdd OAI22X1
X71 NOR2X1_3/Y INVX1_4/gnd NOR2X1_3/A NOR2X1_3/B INVX1_4/vdd NOR2X1
X72 INVX1_5/Y INVX1_4/gnd INVX1_5/A INVX1_4/vdd INVX1
X73 AOI22X1_3/A INVX1_4/gnd INVX1_1/Y INVX1_4/Y OR2X1_1/B INVX1_4/vdd OAI21X1
X74 OR2X1_4/Y INVX1_4/gnd INVX1_4/A OR2X1_4/B INVX1_4/vdd OR2X1
X75 INVX1_4/Y INVX1_4/gnd INVX1_4/A INVX1_4/vdd INVX1
X76 NOR2X1_3/B INVX1_4/gnd INVX1_25/Y INVX1_4/A INVX1_4/vdd NAND2X1
X77 INVX1_25/Y INVX1_4/gnd OR2X1_4/B INVX1_4/vdd INVX1
X78 INVX1_4/gnd clock OAI22X1_10/Y INVX1_6/A INVX1_2/vdd DFFPOSX1
X79 OAI22X1_10/Y INVX1_4/gnd OAI22X1_3/A INVX1_21/Y INVX1_6/Y OR2X1_1/Y INVX1_2/vdd OAI22X1
X80 OAI22X1_2/Y INVX1_4/gnd INVX1_6/Y OAI22X1_3/A INVX1_8/Y OR2X1_1/Y INVX1_2/vdd OAI22X1
X81 INVX1_21/Y INVX1_4/gnd INVX1_21/A INVX1_2/vdd INVX1
X82 OAI22X1_6/Y INVX1_4/gnd MUX2X1_2/Y OAI22X1_3/A OR2X1_1/Y INVX1_21/Y INVX1_2/vdd OAI22X1
X83 OAI22X1_7/Y INVX1_4/gnd OAI22X1_3/A INVX1_8/Y OR2X1_1/Y INVX1_27/Y INVX1_2/vdd OAI22X1
X84 OR2X1_3/Y INVX1_4/gnd OR2X1_1/B OR2X1_2/Y INVX1_2/vdd OR2X1
X85 MUX2X1_2/Y INVX1_4/gnd INVX1_27/A INVX1_27/Y INVX1_2/vdd MUX2X1_1/Y MUX2X1
X86 INVX1_4/gnd clock OAI22X1_11/Y INVX1_10/A INVX1_2/vdd DFFPOSX1
X87 AOI21X1_4/C INVX1_4/gnd MUX2X1_3/Y INVX1_18/A OR2X1_1/B INVX1_31/Y INVX1_2/vdd OAI22X1
X88 INVX1_31/Y INVX1_4/gnd INVX1_31/A INVX1_2/vdd INVX1
X89 INVX1_32/A INVX1_4/gnd INVX1_1/A NOR2X1_2/B AOI21X1_4/C INVX1_2/vdd AOI21X1
X90 NOR2X1_2/B INVX1_4/gnd INVX1_31/A OAI21X1_7/B OAI21X1_7/C INVX1_2/vdd OAI21X1
X91 OAI21X1_7/C INVX1_4/gnd OAI21X1_7/B INVX1_31/A INVX1_2/vdd NAND2X1
X92 INVX1_4/gnd clock OAI21X1_4/Y OR2X1_5/A INVX1_2/vdd DFFPOSX1
X93 INVX1_33/A INVX1_4/gnd INVX1_1/A NOR2X1_4/B AOI21X1_5/C INVX1_2/vdd AOI21X1
X94 INVX1_18/A INVX1_4/gnd INVX1_1/Y OR2X1_1/B INVX1_2/vdd NAND2X1
X95 INVX1_20/Y INVX1_4/gnd INVX1_20/A INVX1_2/vdd INVX1
X96 AOI21X1_5/C INVX1_4/gnd OR2X1_1/B INVX1_20/Y NAND3X1_7/Y INVX1_2/vdd OAI21X1
X97 NOR2X1_4/B INVX1_4/gnd OR2X1_5/B NAND2X1_17/Y INVX1_2/vdd NAND2X1
X98 OR2X1_5/B INVX1_4/gnd NOR2X1_1/Y INVX1_19/Y INVX1_20/Y INVX1_2/vdd NAND3X1
X99 AOI21X1_7/C INVX1_4/gnd AOI22X1_5/Y INVX1_18/A OR2X1_1/B INVX1_38/Y INVX1_2/vdd OAI22X1
X100 INVX1_38/Y INVX1_4/gnd OR2X1_6/A INVX1_2/vdd INVX1
X101 OR2X1_6/B INVX1_4/gnd INVX1_19/Y NOR2X1_3/A INVX1_2/vdd NAND2X1
X102 NOR2X1_1/Y INVX1_4/gnd OR2X1_6/A OR2X1_4/Y INVX1_2/vdd NOR2X1
X103 OAI21X1_17/Y INVX1_4/gnd INVX1_1/Y OR2X1_4/Y AOI22X1_3/Y INVX1_2/vdd OAI21X1
X104 AOI22X1_3/Y INVX1_4/gnd AOI22X1_3/A OR2X1_4/B AOI22X1_3/C INVX1_18/Y INVX1_2/vdd AOI22X1
X105 INVX1_4/gnd clock OAI21X1_17/Y OR2X1_4/B INVX1_2/vdd DFFPOSX1
X106 dp<1> INVX1_2/gnd BUFX2_1/A INVX1_2/vdd BUFX2
X107 INVX1_2/gnd clock OAI21X1_5/Y BUFX2_1/A INVX1_2/vdd DFFPOSX1
X108 OAI21X1_5/C INVX1_2/gnd OR2X1_2/Y BUFX2_1/A INVX1_2/vdd NAND2X1
X109 OAI21X1_5/Y INVX1_2/gnd OR2X1_3/Y INVX1_21/Y OAI21X1_5/C INVX1_2/vdd OAI21X1
X110 INVX1_2/gnd clock OAI22X1_2/Y INVX1_8/A INVX1_2/vdd DFFPOSX1
X111 INVX1_8/Y INVX1_2/gnd INVX1_8/A INVX1_2/vdd INVX1
X112 OAI21X1_10/Y INVX1_2/gnd OR2X1_3/Y INVX1_27/Y OAI21X1_10/C INVX1_2/vdd OAI21X1
X113 OAI21X1_21/Y INVX1_2/gnd INVX1_8/Y OR2X1_3/Y NAND2X1_25/Y INVX1_2/vdd OAI21X1
X114 NAND2X1_25/Y INVX1_2/gnd OR2X1_2/Y BUFX2_2/A INVX1_2/vdd NAND2X1
X115 MUX2X1_3/B INVX1_2/gnd N<8> INVX1_2/vdd INVX1
X116 MUX2X1_3/Y INVX1_2/gnd MUX2X1_3/B N<8> INVX1_2/vdd MUX2X1_3/S MUX2X1
X117 INVX1_22/Y INVX1_2/gnd INVX1_22/A INVX1_2/vdd INVX1
X118 OAI21X1_7/B INVX1_2/gnd INVX1_22/Y NOR2X1_2/A INVX1_2/vdd NAND2X1
X119 AOI21X1_6/C INVX1_2/gnd AOI22X1_4/Y INVX1_18/A OR2X1_1/B INVX1_22/Y INVX1_2/vdd OAI22X1
X120 INVX1_36/A INVX1_2/gnd INVX1_1/A NOR2X1_2/A AOI21X1_6/C INVX1_2/vdd AOI21X1
X121 NOR2X1_2/Y INVX1_2/gnd NOR2X1_2/A NOR2X1_2/B INVX1_2/vdd NOR2X1
X122 NOR2X1_2/A INVX1_2/gnd INVX1_22/A OR2X1_5/Y NAND2X1_9/Y INVX1_2/vdd OAI21X1
X123 NAND2X1_9/Y INVX1_2/gnd OR2X1_5/Y INVX1_22/A INVX1_2/vdd NAND2X1
X124 INVX1_24/A INVX1_2/gnd NOR2X1_2/Y OR2X1_1/B INVX1_23/Y INVX1_2/vdd NAND3X1
X125 INVX1_23/Y INVX1_2/gnd INVX1_23/A INVX1_2/vdd INVX1
X126 OAI21X1_4/Y INVX1_2/gnd OR2X1_1/B INVX1_11/Y AOI22X1_1/Y INVX1_2/vdd OAI21X1
X127 AOI22X1_1/Y INVX1_2/gnd AOI22X1_1/A INVX1_18/Y INVX1_1/A INVX1_23/A INVX1_2/vdd AOI22X1
X128 INVX1_23/A INVX1_2/gnd OR2X1_5/Y NAND2X1_6/Y INVX1_2/vdd NAND2X1
X129 NAND3X1_7/Y INVX1_2/gnd NAND3X1_7/A OR2X1_7/B INVX1_18/Y INVX1_2/vdd NAND3X1
X130 INVX1_11/Y INVX1_2/gnd OR2X1_5/A INVX1_2/vdd INVX1
X131 OR2X1_5/Y INVX1_2/gnd OR2X1_5/A OR2X1_5/B INVX1_2/vdd OR2X1
X132 NAND2X1_6/Y INVX1_2/gnd OR2X1_5/B OR2X1_5/A INVX1_2/vdd NAND2X1
X133 INVX1_18/Y INVX1_2/gnd INVX1_18/A INVX1_2/vdd INVX1
X134 INVX1_26/A INVX1_2/gnd INVX1_1/A NOR2X1_3/A AOI21X1_3/C INVX1_2/vdd AOI21X1
X135 AOI21X1_3/C INVX1_2/gnd OAI22X1_5/A INVX1_18/A OR2X1_1/B INVX1_19/Y INVX1_2/vdd OAI22X1
X136 INVX1_19/Y INVX1_2/gnd INVX1_19/A INVX1_2/vdd INVX1
X137 NOR2X1_3/A INVX1_2/gnd INVX1_19/A OR2X1_4/Y OAI21X1_8/C INVX1_2/vdd OAI21X1
X138 OAI21X1_8/C INVX1_2/gnd OR2X1_4/Y INVX1_19/A INVX1_2/vdd NAND2X1
X139 INVX1_2/Y INVX1_2/gnd N<1> INVX1_2/vdd INVX1
X140 AOI22X1_3/C INVX1_2/gnd N<1> N<2> NOR2X1_5/B INVX1_2/vdd OAI21X1
X141 NOR2X1_5/B INVX1_2/gnd N<1> N<2> INVX1_2/vdd NAND2X1
X142 dp<0> INVX1_2/gnd BUFX2_6/A OR2X1_7/vdd BUFX2
X143 INVX1_2/gnd clock OAI21X1_20/Y BUFX2_6/A OR2X1_7/vdd DFFPOSX1
X144 OAI21X1_20/C INVX1_2/gnd OR2X1_2/Y BUFX2_6/A OR2X1_7/vdd NAND2X1
X145 OAI21X1_20/Y INVX1_2/gnd OR2X1_2/Y INVX1_37/Y OAI21X1_20/C OR2X1_7/vdd OAI21X1
X146 INVX1_37/Y INVX1_2/gnd N<0> OR2X1_7/vdd INVX1
X147 dp<4> INVX1_2/gnd BUFX2_8/A OR2X1_7/vdd BUFX2
X148 INVX1_2/gnd clock OAI21X1_10/Y BUFX2_8/A OR2X1_7/vdd DFFPOSX1
X149 OAI21X1_10/C INVX1_2/gnd OR2X1_2/Y BUFX2_8/A OR2X1_7/vdd NAND2X1
X150 INVX1_2/gnd clock OAI21X1_21/Y BUFX2_2/A OR2X1_7/vdd DFFPOSX1
X151 dp<3> INVX1_2/gnd BUFX2_2/A OR2X1_7/vdd BUFX2
X152 MUX2X1_3/S INVX1_2/gnd N<7> OR2X1_7/Y OR2X1_7/vdd NOR2X1
X153 AOI22X1_4/Y INVX1_2/gnd N<7> INVX1_34/Y INVX1_35/Y OR2X1_7/Y OR2X1_7/vdd AOI22X1
X154 INVX1_35/Y INVX1_2/gnd N<7> OR2X1_7/vdd INVX1
X155 INVX1_34/Y INVX1_2/gnd OR2X1_7/Y OR2X1_7/vdd INVX1
X156 INVX1_36/Y INVX1_2/gnd INVX1_36/A OR2X1_7/vdd INVX1
X157 INVX1_2/gnd clock INVX1_36/Y INVX1_22/A OR2X1_7/vdd DFFPOSX1
X158 OR2X1_7/Y INVX1_2/gnd N<6> OR2X1_7/B OR2X1_7/vdd OR2X1
X159 INVX1_17/Y INVX1_2/gnd N<6> OR2X1_7/vdd INVX1
X160 AOI22X1_1/A INVX1_2/gnd N<6> INVX1_16/Y INVX1_17/Y OR2X1_7/B OR2X1_7/vdd OAI22X1
X161 INVX1_16/Y INVX1_2/gnd OR2X1_7/B OR2X1_7/vdd INVX1
X162 INVX1_15/Y INVX1_2/gnd N<5> OR2X1_7/vdd INVX1
X163 OR2X1_7/B INVX1_2/gnd INVX1_13/Y INVX1_14/Y INVX1_15/Y OR2X1_7/vdd NAND3X1
X164 INVX1_14/Y INVX1_2/gnd N<4> OR2X1_7/vdd INVX1
X165 NAND3X1_7/A INVX1_2/gnd N<4> INVX1_13/A N<5> OR2X1_7/vdd OAI21X1
X166 INVX1_13/Y INVX1_2/gnd INVX1_13/A OR2X1_7/vdd INVX1
X167 AOI22X1_5/Y INVX1_2/gnd INVX1_13/Y N<4> INVX1_14/Y INVX1_13/A OR2X1_7/vdd AOI22X1
X168 INVX1_26/Y INVX1_2/gnd INVX1_26/A OR2X1_7/vdd INVX1
X169 INVX1_2/gnd clock INVX1_26/Y INVX1_19/A OR2X1_7/vdd DFFPOSX1
X170 INVX1_13/A INVX1_2/gnd INVX1_12/Y NOR2X1_5/B OR2X1_7/vdd NAND2X1
X171 INVX1_12/Y INVX1_2/gnd N<3> OR2X1_7/vdd INVX1
X172 OAI22X1_5/A INVX1_2/gnd NOR2X1_5/B N<3> NOR2X1_5/Y OR2X1_7/vdd AOI21X1
X173 NOR2X1_5/Y INVX1_2/gnd N<3> NOR2X1_5/B OR2X1_7/vdd NOR2X1
.end

