* hier1.spice--- with hier2.spice, mixed-hierarchy LVS test

.subckt invert in1 out1 Vdd Gnd
M1 out1 in1 Vdd Vdd pmos w=800n l=400n
M2 out1 in1 Gnd Gnd nmos w=800n l=400n
.ends

.subckt buffer in1 out1 Vdd Gnd
X1 in1 mid Vdd Gnd invert
X2 mid out1 Vdd Gnd invert
.ends

X1 in out Vdd Gnd buffer

